V1 1 0 dc 20
R1 1 2 5k
R2 2 0 4k
R3 3 0 1k
I1 3 2 2mA
.op
.end
